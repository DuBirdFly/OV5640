module shift_custom (
    input  wire                         vga_clk                    ,
    input  wire                         rst_n                      ,
    ports
);


























endmodule
